`default_nettype none
`timescale 1ns/1ps

`ifndef RIP_COMMON
`define RIP_COMMON

package rip_common;
    `include "rip_const.svh"
    `include "rip_type.svh"
endpackage: rip_common

`endif  // RIP_COMMON
